-------------------------------------------
-- Delivery #21
-- Fabrício da Costa Guimarães - 21950515
-- Perfil Comportamental: LOBO
-- Engenharia da Computação - FT UFAM
-- ED2 e LED - 2021/01 - Equipe 06
-------------------------------------------

-- Bibliotecas e pacotes
use work.dsf_std.all;

-- Entidade
entity logic_h0 is
	port(
		gt: in bit; 
		lt: in bit; 
	
		q: buffer bit
	);
end entity logic_h0;

-- Arquitetura
architecture logic_h0_a of logic_h0 is
begin
-- vazia
	
end architecture logic_h0_a;